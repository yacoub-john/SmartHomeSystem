pll_ip	pll_inst (
	.inclk0 ( inclk0_sig ),
	.c0 ( c0_sig ),
	.c1 ( c1_sig ),
	.c2 ( c2_sig )
	);
